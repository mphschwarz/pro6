module AC_MOTOR_SINE_SECTOR(
	input CLK,
	input [bits - 1:0] FREQUENCY,
	output reg [2:0] SECTOR,
	output reg [bits - 1:0] SINE_POSITIVE,
	output reg [bits - 1:0] SINE_NEGATIVE
);

parameter sine_samples = 512 * 6;
parameter bits = 12;

parameter f_clk = 100 * 10**6;
parameter f_min = 12;
parameter f_max = 60;
parameter clock_div_min =  f_clk / (f_min * sine_samples);
parameter clock_div_max =  f_clk / (f_max * sine_samples);

reg [12:0] clock_div;
reg [8:0] memory_pos;
reg [8:0] memory_neg;
reg [12:0] freq_int;

(* ramstyle = "M9K" *) reg [bits-1:0] sine [(sine_samples / 6) - 1:0];

always @(posedge CLK) begin
	freq_int <= FREQUENCY + clock_div_max;
end

always @(posedge CLK) begin
	if (clock_div >= freq_int) begin // increment RAM-pointers
		clock_div <= 0;
		memory_pos <= memory_pos + 1;
		memory_neg <= memory_neg - 1;
	end else begin
		clock_div <= clock_div + 1;
	end
end

always @(posedge CLK) begin
	// increment sector at last clock cycle
	if(memory_pos == 0/*sine_samples / 6 - 1*/ && clock_div == 0 /*freq_int*/) begin
		if (SECTOR == 5) begin
			SECTOR <= 0;
		end else begin 
			SECTOR <= SECTOR + 1;
		end
	end
end

always @(posedge CLK) begin
	SINE_POSITIVE <= sine[memory_pos];
	SINE_NEGATIVE <= sine[memory_neg];
end

initial begin
	clock_div <= 0;
	memory_pos <= 0;
	memory_neg <= 2**9 - 1;
	freq_int <= 0;
	SECTOR <= 0;
	SINE_POSITIVE <= 0;
	SINE_NEGATIVE <= 12'b110111011000;

	sine[0] = 12'b000000000100; sine[1] = 12'b000000001100;
	sine[2] = 12'b000000010100; sine[3] = 12'b000000011101;
	sine[4] = 12'b000000100101; sine[5] = 12'b000000101110;
	sine[6] = 12'b000000110110; sine[7] = 12'b000000111110;
	sine[8] = 12'b000001000111; sine[9] = 12'b000001001111;
	sine[10] = 12'b000001010111; sine[11] = 12'b000001100000;
	sine[12] = 12'b000001101000; sine[13] = 12'b000001110001;
	sine[14] = 12'b000001111001; sine[15] = 12'b000010000001;
	sine[16] = 12'b000010001010; sine[17] = 12'b000010010010;
	sine[18] = 12'b000010011010; sine[19] = 12'b000010100011;
	sine[20] = 12'b000010101011; sine[21] = 12'b000010110100;
	sine[22] = 12'b000010111100; sine[23] = 12'b000011000100;
	sine[24] = 12'b000011001101; sine[25] = 12'b000011010101;
	sine[26] = 12'b000011011101; sine[27] = 12'b000011100110;
	sine[28] = 12'b000011101110; sine[29] = 12'b000011110110;
	sine[30] = 12'b000011111111; sine[31] = 12'b000100000111;
	sine[32] = 12'b000100010000; sine[33] = 12'b000100011000;
	sine[34] = 12'b000100100000; sine[35] = 12'b000100101001;
	sine[36] = 12'b000100110001; sine[37] = 12'b000100111001;
	sine[38] = 12'b000101000010; sine[39] = 12'b000101001010;
	sine[40] = 12'b000101010010; sine[41] = 12'b000101011011;
	sine[42] = 12'b000101100011; sine[43] = 12'b000101101011;
	sine[44] = 12'b000101110100; sine[45] = 12'b000101111100;
	sine[46] = 12'b000110000100; sine[47] = 12'b000110001101;
	sine[48] = 12'b000110010101; sine[49] = 12'b000110011101;
	sine[50] = 12'b000110100110; sine[51] = 12'b000110101110;
	sine[52] = 12'b000110110110; sine[53] = 12'b000110111111;
	sine[54] = 12'b000111000111; sine[55] = 12'b000111001111;
	sine[56] = 12'b000111011000; sine[57] = 12'b000111100000;
	sine[58] = 12'b000111101000; sine[59] = 12'b000111110001;
	sine[60] = 12'b000111111001; sine[61] = 12'b001000000001;
	sine[62] = 12'b001000001010; sine[63] = 12'b001000010010;
	sine[64] = 12'b001000011010; sine[65] = 12'b001000100010;
	sine[66] = 12'b001000101011; sine[67] = 12'b001000110011;
	sine[68] = 12'b001000111011; sine[69] = 12'b001001000100;
	sine[70] = 12'b001001001100; sine[71] = 12'b001001010100;
	sine[72] = 12'b001001011101; sine[73] = 12'b001001100101;
	sine[74] = 12'b001001101101; sine[75] = 12'b001001110101;
	sine[76] = 12'b001001111110; sine[77] = 12'b001010000110;
	sine[78] = 12'b001010001110; sine[79] = 12'b001010010110;
	sine[80] = 12'b001010011111; sine[81] = 12'b001010100111;
	sine[82] = 12'b001010101111; sine[83] = 12'b001010110111;
	sine[84] = 12'b001011000000; sine[85] = 12'b001011001000;
	sine[86] = 12'b001011010000; sine[87] = 12'b001011011000;
	sine[88] = 12'b001011100001; sine[89] = 12'b001011101001;
	sine[90] = 12'b001011110001; sine[91] = 12'b001011111001;
	sine[92] = 12'b001100000010; sine[93] = 12'b001100001010;
	sine[94] = 12'b001100010010; sine[95] = 12'b001100011010;
	sine[96] = 12'b001100100011; sine[97] = 12'b001100101011;
	sine[98] = 12'b001100110011; sine[99] = 12'b001100111011;
	sine[100] = 12'b001101000011; sine[101] = 12'b001101001100;
	sine[102] = 12'b001101010100; sine[103] = 12'b001101011100;
	sine[104] = 12'b001101100100; sine[105] = 12'b001101101100;
	sine[106] = 12'b001101110100; sine[107] = 12'b001101111101;
	sine[108] = 12'b001110000101; sine[109] = 12'b001110001101;
	sine[110] = 12'b001110010101; sine[111] = 12'b001110011101;
	sine[112] = 12'b001110100101; sine[113] = 12'b001110101110;
	sine[114] = 12'b001110110110; sine[115] = 12'b001110111110;
	sine[116] = 12'b001111000110; sine[117] = 12'b001111001110;
	sine[118] = 12'b001111010110; sine[119] = 12'b001111011110;
	sine[120] = 12'b001111100111; sine[121] = 12'b001111101111;
	sine[122] = 12'b001111110111; sine[123] = 12'b001111111111;
	sine[124] = 12'b010000000111; sine[125] = 12'b010000001111;
	sine[126] = 12'b010000010111; sine[127] = 12'b010000011111;
	sine[128] = 12'b010000100111; sine[129] = 12'b010000101111;
	sine[130] = 12'b010000111000; sine[131] = 12'b010001000000;
	sine[132] = 12'b010001001000; sine[133] = 12'b010001010000;
	sine[134] = 12'b010001011000; sine[135] = 12'b010001100000;
	sine[136] = 12'b010001101000; sine[137] = 12'b010001110000;
	sine[138] = 12'b010001111000; sine[139] = 12'b010010000000;
	sine[140] = 12'b010010001000; sine[141] = 12'b010010010000;
	sine[142] = 12'b010010011000; sine[143] = 12'b010010100000;
	sine[144] = 12'b010010101000; sine[145] = 12'b010010110000;
	sine[146] = 12'b010010111000; sine[147] = 12'b010011000000;
	sine[148] = 12'b010011001000; sine[149] = 12'b010011010000;
	sine[150] = 12'b010011011000; sine[151] = 12'b010011100000;
	sine[152] = 12'b010011101000; sine[153] = 12'b010011110000;
	sine[154] = 12'b010011111000; sine[155] = 12'b010100000000;
	sine[156] = 12'b010100001000; sine[157] = 12'b010100010000;
	sine[158] = 12'b010100011000; sine[159] = 12'b010100100000;
	sine[160] = 12'b010100101000; sine[161] = 12'b010100110000;
	sine[162] = 12'b010100111000; sine[163] = 12'b010101000000;
	sine[164] = 12'b010101000111; sine[165] = 12'b010101001111;
	sine[166] = 12'b010101010111; sine[167] = 12'b010101011111;
	sine[168] = 12'b010101100111; sine[169] = 12'b010101101111;
	sine[170] = 12'b010101110111; sine[171] = 12'b010101111111;
	sine[172] = 12'b010110000110; sine[173] = 12'b010110001110;
	sine[174] = 12'b010110010110; sine[175] = 12'b010110011110;
	sine[176] = 12'b010110100110; sine[177] = 12'b010110101110;
	sine[178] = 12'b010110110110; sine[179] = 12'b010110111101;
	sine[180] = 12'b010111000101; sine[181] = 12'b010111001101;
	sine[182] = 12'b010111010101; sine[183] = 12'b010111011101;
	sine[184] = 12'b010111100100; sine[185] = 12'b010111101100;
	sine[186] = 12'b010111110100; sine[187] = 12'b010111111100;
	sine[188] = 12'b011000000011; sine[189] = 12'b011000001011;
	sine[190] = 12'b011000010011; sine[191] = 12'b011000011011;
	sine[192] = 12'b011000100010; sine[193] = 12'b011000101010;
	sine[194] = 12'b011000110010; sine[195] = 12'b011000111010;
	sine[196] = 12'b011001000001; sine[197] = 12'b011001001001;
	sine[198] = 12'b011001010001; sine[199] = 12'b011001011000;
	sine[200] = 12'b011001100000; sine[201] = 12'b011001101000;
	sine[202] = 12'b011001101111; sine[203] = 12'b011001110111;
	sine[204] = 12'b011001111111; sine[205] = 12'b011010000110;
	sine[206] = 12'b011010001110; sine[207] = 12'b011010010110;
	sine[208] = 12'b011010011101; sine[209] = 12'b011010100101;
	sine[210] = 12'b011010101101; sine[211] = 12'b011010110100;
	sine[212] = 12'b011010111100; sine[213] = 12'b011011000011;
	sine[214] = 12'b011011001011; sine[215] = 12'b011011010011;
	sine[216] = 12'b011011011010; sine[217] = 12'b011011100010;
	sine[218] = 12'b011011101001; sine[219] = 12'b011011110001;
	sine[220] = 12'b011011111000; sine[221] = 12'b011100000000;
	sine[222] = 12'b011100000111; sine[223] = 12'b011100001111;
	sine[224] = 12'b011100010110; sine[225] = 12'b011100011110;
	sine[226] = 12'b011100100101; sine[227] = 12'b011100101101;
	sine[228] = 12'b011100110100; sine[229] = 12'b011100111100;
	sine[230] = 12'b011101000011; sine[231] = 12'b011101001011;
	sine[232] = 12'b011101010010; sine[233] = 12'b011101011010;
	sine[234] = 12'b011101100001; sine[235] = 12'b011101101001;
	sine[236] = 12'b011101110000; sine[237] = 12'b011101110111;
	sine[238] = 12'b011101111111; sine[239] = 12'b011110000110;
	sine[240] = 12'b011110001110; sine[241] = 12'b011110010101;
	sine[242] = 12'b011110011100; sine[243] = 12'b011110100100;
	sine[244] = 12'b011110101011; sine[245] = 12'b011110110010;
	sine[246] = 12'b011110111010; sine[247] = 12'b011111000001;
	sine[248] = 12'b011111001000; sine[249] = 12'b011111010000;
	sine[250] = 12'b011111010111; sine[251] = 12'b011111011110;
	sine[252] = 12'b011111100110; sine[253] = 12'b011111101101;
	sine[254] = 12'b011111110100; sine[255] = 12'b011111111011;
	sine[256] = 12'b100000000011; sine[257] = 12'b100000001010;
	sine[258] = 12'b100000010001; sine[259] = 12'b100000011000;
	sine[260] = 12'b100000100000; sine[261] = 12'b100000100111;
	sine[262] = 12'b100000101110; sine[263] = 12'b100000110101;
	sine[264] = 12'b100000111100; sine[265] = 12'b100001000100;
	sine[266] = 12'b100001001011; sine[267] = 12'b100001010010;
	sine[268] = 12'b100001011001; sine[269] = 12'b100001100000;
	sine[270] = 12'b100001100111; sine[271] = 12'b100001101110;
	sine[272] = 12'b100001110101; sine[273] = 12'b100001111101;
	sine[274] = 12'b100010000100; sine[275] = 12'b100010001011;
	sine[276] = 12'b100010010010; sine[277] = 12'b100010011001;
	sine[278] = 12'b100010100000; sine[279] = 12'b100010100111;
	sine[280] = 12'b100010101110; sine[281] = 12'b100010110101;
	sine[282] = 12'b100010111100; sine[283] = 12'b100011000011;
	sine[284] = 12'b100011001010; sine[285] = 12'b100011010001;
	sine[286] = 12'b100011011000; sine[287] = 12'b100011011111;
	sine[288] = 12'b100011100110; sine[289] = 12'b100011101101;
	sine[290] = 12'b100011110100; sine[291] = 12'b100011111011;
	sine[292] = 12'b100100000010; sine[293] = 12'b100100001001;
	sine[294] = 12'b100100010000; sine[295] = 12'b100100010111;
	sine[296] = 12'b100100011101; sine[297] = 12'b100100100100;
	sine[298] = 12'b100100101011; sine[299] = 12'b100100110010;
	sine[300] = 12'b100100111001; sine[301] = 12'b100101000000;
	sine[302] = 12'b100101000111; sine[303] = 12'b100101001101;
	sine[304] = 12'b100101010100; sine[305] = 12'b100101011011;
	sine[306] = 12'b100101100010; sine[307] = 12'b100101101001;
	sine[308] = 12'b100101101111; sine[309] = 12'b100101110110;
	sine[310] = 12'b100101111101; sine[311] = 12'b100110000100;
	sine[312] = 12'b100110001010; sine[313] = 12'b100110010001;
	sine[314] = 12'b100110011000; sine[315] = 12'b100110011110;
	sine[316] = 12'b100110100101; sine[317] = 12'b100110101100;
	sine[318] = 12'b100110110010; sine[319] = 12'b100110111001;
	sine[320] = 12'b100111000000; sine[321] = 12'b100111000110;
	sine[322] = 12'b100111001101; sine[323] = 12'b100111010100;
	sine[324] = 12'b100111011010; sine[325] = 12'b100111100001;
	sine[326] = 12'b100111100111; sine[327] = 12'b100111101110;
	sine[328] = 12'b100111110100; sine[329] = 12'b100111111011;
	sine[330] = 12'b101000000010; sine[331] = 12'b101000001000;
	sine[332] = 12'b101000001111; sine[333] = 12'b101000010101;
	sine[334] = 12'b101000011100; sine[335] = 12'b101000100010;
	sine[336] = 12'b101000101001; sine[337] = 12'b101000101111;
	sine[338] = 12'b101000110101; sine[339] = 12'b101000111100;
	sine[340] = 12'b101001000010; sine[341] = 12'b101001001001;
	sine[342] = 12'b101001001111; sine[343] = 12'b101001010110;
	sine[344] = 12'b101001011100; sine[345] = 12'b101001100010;
	sine[346] = 12'b101001101001; sine[347] = 12'b101001101111;
	sine[348] = 12'b101001110101; sine[349] = 12'b101001111100;
	sine[350] = 12'b101010000010; sine[351] = 12'b101010001000;
	sine[352] = 12'b101010001111; sine[353] = 12'b101010010101;
	sine[354] = 12'b101010011011; sine[355] = 12'b101010100001;
	sine[356] = 12'b101010101000; sine[357] = 12'b101010101110;
	sine[358] = 12'b101010110100; sine[359] = 12'b101010111010;
	sine[360] = 12'b101011000001; sine[361] = 12'b101011000111;
	sine[362] = 12'b101011001101; sine[363] = 12'b101011010011;
	sine[364] = 12'b101011011001; sine[365] = 12'b101011011111;
	sine[366] = 12'b101011100110; sine[367] = 12'b101011101100;
	sine[368] = 12'b101011110010; sine[369] = 12'b101011111000;
	sine[370] = 12'b101011111110; sine[371] = 12'b101100000100;
	sine[372] = 12'b101100001010; sine[373] = 12'b101100010000;
	sine[374] = 12'b101100010110; sine[375] = 12'b101100011100;
	sine[376] = 12'b101100100010; sine[377] = 12'b101100101000;
	sine[378] = 12'b101100101110; sine[379] = 12'b101100110100;
	sine[380] = 12'b101100111010; sine[381] = 12'b101101000000;
	sine[382] = 12'b101101000110; sine[383] = 12'b101101001100;
	sine[384] = 12'b101101010010; sine[385] = 12'b101101011000;
	sine[386] = 12'b101101011110; sine[387] = 12'b101101100100;
	sine[388] = 12'b101101101010; sine[389] = 12'b101101101111;
	sine[390] = 12'b101101110101; sine[391] = 12'b101101111011;
	sine[392] = 12'b101110000001; sine[393] = 12'b101110000111;
	sine[394] = 12'b101110001101; sine[395] = 12'b101110010010;
	sine[396] = 12'b101110011000; sine[397] = 12'b101110011110;
	sine[398] = 12'b101110100100; sine[399] = 12'b101110101001;
	sine[400] = 12'b101110101111; sine[401] = 12'b101110110101;
	sine[402] = 12'b101110111011; sine[403] = 12'b101111000000;
	sine[404] = 12'b101111000110; sine[405] = 12'b101111001100;
	sine[406] = 12'b101111010001; sine[407] = 12'b101111010111;
	sine[408] = 12'b101111011101; sine[409] = 12'b101111100010;
	sine[410] = 12'b101111101000; sine[411] = 12'b101111101101;
	sine[412] = 12'b101111110011; sine[413] = 12'b101111111000;
	sine[414] = 12'b101111111110; sine[415] = 12'b110000000100;
	sine[416] = 12'b110000001001; sine[417] = 12'b110000001111;
	sine[418] = 12'b110000010100; sine[419] = 12'b110000011010;
	sine[420] = 12'b110000011111; sine[421] = 12'b110000100100;
	sine[422] = 12'b110000101010; sine[423] = 12'b110000101111;
	sine[424] = 12'b110000110101; sine[425] = 12'b110000111010;
	sine[426] = 12'b110001000000; sine[427] = 12'b110001000101;
	sine[428] = 12'b110001001010; sine[429] = 12'b110001010000;
	sine[430] = 12'b110001010101; sine[431] = 12'b110001011010;
	sine[432] = 12'b110001100000; sine[433] = 12'b110001100101;
	sine[434] = 12'b110001101010; sine[435] = 12'b110001101111;
	sine[436] = 12'b110001110101; sine[437] = 12'b110001111010;
	sine[438] = 12'b110001111111; sine[439] = 12'b110010000100;
	sine[440] = 12'b110010001010; sine[441] = 12'b110010001111;
	sine[442] = 12'b110010010100; sine[443] = 12'b110010011001;
	sine[444] = 12'b110010011110; sine[445] = 12'b110010100011;
	sine[446] = 12'b110010101001; sine[447] = 12'b110010101110;
	sine[448] = 12'b110010110011; sine[449] = 12'b110010111000;
	sine[450] = 12'b110010111101; sine[451] = 12'b110011000010;
	sine[452] = 12'b110011000111; sine[453] = 12'b110011001100;
	sine[454] = 12'b110011010001; sine[455] = 12'b110011010110;
	sine[456] = 12'b110011011011; sine[457] = 12'b110011100000;
	sine[458] = 12'b110011100101; sine[459] = 12'b110011101010;
	sine[460] = 12'b110011101111; sine[461] = 12'b110011110100;
	sine[462] = 12'b110011111001; sine[463] = 12'b110011111110;
	sine[464] = 12'b110100000011; sine[465] = 12'b110100000111;
	sine[466] = 12'b110100001100; sine[467] = 12'b110100010001;
	sine[468] = 12'b110100010110; sine[469] = 12'b110100011011;
	sine[470] = 12'b110100100000; sine[471] = 12'b110100100100;
	sine[472] = 12'b110100101001; sine[473] = 12'b110100101110;
	sine[474] = 12'b110100110011; sine[475] = 12'b110100110111;
	sine[476] = 12'b110100111100; sine[477] = 12'b110101000001;
	sine[478] = 12'b110101000101; sine[479] = 12'b110101001010;
	sine[480] = 12'b110101001111; sine[481] = 12'b110101010011;
	sine[482] = 12'b110101011000; sine[483] = 12'b110101011101;
	sine[484] = 12'b110101100001; sine[485] = 12'b110101100110;
	sine[486] = 12'b110101101010; sine[487] = 12'b110101101111;
	sine[488] = 12'b110101110011; sine[489] = 12'b110101111000;
	sine[490] = 12'b110101111100; sine[491] = 12'b110110000001;
	sine[492] = 12'b110110000101; sine[493] = 12'b110110001010;
	sine[494] = 12'b110110001110; sine[495] = 12'b110110010011;
	sine[496] = 12'b110110010111; sine[497] = 12'b110110011100;
	sine[498] = 12'b110110100000; sine[499] = 12'b110110100100;
	sine[500] = 12'b110110101001; sine[501] = 12'b110110101101;
	sine[502] = 12'b110110110001; sine[503] = 12'b110110110110;
	sine[504] = 12'b110110111010; sine[505] = 12'b110110111110;
	sine[506] = 12'b110111000011; sine[507] = 12'b110111000111;
	sine[508] = 12'b110111001011; sine[509] = 12'b110111001111;
	sine[510] = 12'b110111010100; sine[511] = 12'b110111011000;
	
end
endmodule
