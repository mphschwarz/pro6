////////////////////////////////////////////////////////////////////////////////////////////
module MAX_12_BIT(
	input CLK,
	input [11:0] IN_1,
	input [11:0] IN_2,
	output reg [11:0] OUT);
	//
	initial
		begin
			OUT <= 0;
		end
	//
	always @(posedge CLK)
	begin	
		if (IN_1 >= IN_2) OUT <= IN_1;
		else OUT <= IN_2;
	end
endmodule
////////////////////////////////////////////////////////////////////////////////////////////