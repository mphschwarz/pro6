module AC_MOTOR_MODULAR(
	input CLK,
	input ENABLE,
	
	input CW,
	input CCW,
	input FREQUENCY,
	input AMPLITUDE,

	output OUT1,
	output OUT2,
	output OUT3,
	output OUT4,
	output OUT5,
	output OUT6,
	
	output EN1,
	output EN2,
	output EN3,
	output EN4,
	output EN5,
	output EN6);

	assign EN1 = 1;
	assign EN2 = 1;
	assign EN3 = 1;
	assign EN4 = 1;
	assign EN5 = 1;
	assign EN6 = 1;


